library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity template is
Port (	clk : in STD_LOGIC;
		rst : in STD_LOGIC
	 );
end template;

architecture Behavioral of template is

begin

end Behavioral;

